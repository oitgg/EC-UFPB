CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 100 9
0 71 1366 728
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1366 728
143654930 0
0
6 Title:
5 Name:
0
0
0
22
8 3-In OR~
219 534 456 0 4 22
0 11 10 9 8
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 7 0
1 U
8953 0 0
0
0
9 2-In XOR~
219 549 325 0 3 22
0 13 7 12
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 6 0
1 U
4441 0 0
0
0
9 2-In AND~
219 468 505 0 3 22
0 3 2 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 5 0
1 U
3618 0 0
0
0
9 2-In AND~
219 469 461 0 3 22
0 4 3 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 3 0
1 U
6153 0 0
0
0
9 2-In AND~
219 467 418 0 3 22
0 4 2 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 3 0
1 U
5394 0 0
0
0
9 Inverter~
13 298 353 0 2 22
0 6 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 2 0
1 U
7734 0 0
0
0
9 2-In XOR~
219 637 330 0 3 22
0 12 8 14
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 1 0
1 U
9914 0 0
0
0
9 2-In XOR~
219 531 229 0 3 22
0 2 17 15
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 1 0
1 U
3747 0 0
0
0
9 2-In AND~
219 412 196 0 3 22
0 18 5 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
3549 0 0
0
0
12 Hex Display~
7 42 490 0 18 19
10 5 3 7 20 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
1 Y
-4 -38 3 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
7931 0 0
0
0
8 Hex Key~
166 132 562 0 11 12
0 7 21 22 23 0 0 0 0 0
0 48
0
0 0 4656 0
0
2 B3
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
3 KPD
9325 0 0
0
0
8 Hex Key~
166 132 502 0 11 12
0 3 5 5 5 0 0 0 0 0
1 49
0
0 0 4656 0
0
2 B2
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
8903 0 0
0
0
8 Hex Key~
166 131 437 0 11 12
0 5 24 25 26 0 0 0 0 0
1 49
0
0 0 4656 0
0
2 B1
-6 -35 8 -27
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
3 KPD
3834 0 0
0
0
9 2-In XOR~
219 387 296 0 3 22
0 6 3 17
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
3363 0 0
0
0
9 Inverter~
13 285 163 0 2 22
0 19 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 2 0
1 U
7668 0 0
0
0
9 2-In XOR~
219 348 132 0 3 22
0 19 5 16
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1446731082
65 0 0 0 4 1 1 0
1 U
4718 0 0
0
0
8 Hex Key~
166 141 206 0 11 12
0 13 27 28 29 0 0 0 0 0
1 49
0
0 0 4656 0
0
2 A3
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
3 KPD
3874 0 0
0
0
8 Hex Key~
166 138 139 0 11 12
0 6 30 31 32 0 0 0 0 0
0 48
0
0 0 4656 0
0
2 A2
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
3 KPD
6671 0 0
0
0
8 Hex Key~
166 136 71 0 11 12
0 19 33 34 35 0 0 0 0 0
1 49
0
0 0 4656 0
0
2 A1
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
3 KPD
3789 0 0
0
0
12 Hex Display~
7 728 102 0 18 19
10 16 15 14 36 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
7 Resulta
-25 -38 24 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
4871 0 0
0
0
12 Hex Display~
7 51 171 0 18 19
10 19 6 13 37 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
1 X
-4 -38 3 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
3750 0 0
0
0
7 Ground~
168 24 586 0 1 3
0 38
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 0 0 0 0
3 GND
8778 0 0
0
0
35
2 0 2 0 0 8192 0 3 0 0 4 3
444 514
438 514
438 427
1 0 3 0 0 8192 0 3 0 0 3 3
444 496
426 496
426 470
2 0 3 0 0 4224 0 4 0 0 15 2
445 470
198 470
2 0 2 0 0 8336 0 5 0 0 27 3
443 427
436 427
436 196
1 0 4 0 0 4096 0 4 0 0 13 3
445 452
354 452
354 409
4 0 5 0 0 0 0 12 0 0 12 2
123 526
123 526
3 0 5 0 0 0 0 12 0 0 12 2
129 526
129 526
2 0 5 0 0 0 0 12 0 0 12 2
135 526
135 526
0 1 6 0 0 4096 0 0 6 34 0 4
363 282
275 282
275 353
283 353
0 3 7 0 0 8192 0 0 10 14 0 4
187 590
187 614
39 614
39 514
0 2 3 0 0 0 0 0 10 15 0 4
153 530
153 541
45 541
45 514
0 1 5 0 0 8192 0 0 10 31 0 4
174 465
174 526
51 526
51 514
1 2 4 0 0 4224 0 5 6 0 0 4
443 409
327 409
327 353
319 353
1 2 7 0 0 12416 0 11 2 0 0 5
141 586
141 590
384 590
384 334
533 334
1 2 3 0 0 0 0 12 14 0 0 6
141 526
141 530
198 530
198 298
371 298
371 305
4 2 8 0 0 8320 0 1 7 0 0 4
567 456
613 456
613 339
621 339
3 3 9 0 0 8320 0 3 1 0 0 4
489 505
513 505
513 465
521 465
3 2 10 0 0 4224 0 4 1 0 0 4
490 461
513 461
513 456
522 456
3 1 11 0 0 8320 0 5 1 0 0 4
488 418
513 418
513 447
521 447
3 1 12 0 0 4224 0 2 7 0 0 4
582 325
613 325
613 321
621 321
0 3 13 0 0 4096 0 0 21 22 0 3
150 255
48 255
48 195
1 1 13 0 0 8320 0 17 2 0 0 3
150 230
150 316
533 316
3 3 14 0 0 8320 0 7 20 0 0 3
670 330
725 330
725 126
3 2 15 0 0 8320 0 8 20 0 0 4
564 229
564 155
731 155
731 126
3 1 16 0 0 4224 0 16 20 0 0 3
381 132
737 132
737 126
3 2 17 0 0 4224 0 14 8 0 0 4
420 296
507 296
507 238
515 238
3 1 2 0 0 0 0 9 8 0 0 4
433 196
507 196
507 220
515 220
2 0 5 0 0 4096 0 9 0 0 31 2
388 205
241 205
2 1 18 0 0 4224 0 15 9 0 0 4
306 163
380 163
380 187
388 187
0 1 19 0 0 8192 0 0 15 35 0 3
212 111
212 163
270 163
1 2 5 0 0 12416 0 13 16 0 0 5
140 461
140 465
241 465
241 141
332 141
0 2 6 0 0 8192 0 0 21 34 0 6
162 178
162 170
72 170
72 203
54 203
54 195
0 1 19 0 0 12288 0 0 21 35 0 6
170 111
170 25
72 25
72 203
60 203
60 195
1 1 6 0 0 8320 0 18 14 0 0 5
147 163
147 178
363 178
363 287
371 287
1 1 19 0 0 8320 0 19 16 0 0 5
145 95
145 111
324 111
324 123
332 123
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3999480 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
