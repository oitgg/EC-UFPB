CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 40 30 100 9
0 71 1366 728
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1366 728
143654930 0
0
6 Title:
5 Name:
0
0
0
22
8 3-In OR~
219 552 376 0 4 22
0 12 11 10 9
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 7 0
1 U
8953 0 0
0
0
9 2-In XOR~
219 389 326 0 3 22
0 3 8 13
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 6 0
1 U
4441 0 0
0
0
9 2-In AND~
219 560 506 0 3 22
0 5 4 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 5 0
1 U
3618 0 0
0
0
9 2-In AND~
219 560 469 0 3 22
0 6 5 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-17 -25 4 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 3 0
1 U
6153 0 0
0
0
9 2-In AND~
219 560 426 0 3 22
0 6 4 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 3 0
1 U
5394 0 0
0
0
9 Inverter~
13 298 353 0 2 22
0 7 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 2 0
1 U
7734 0 0
0
0
9 2-In XOR~
219 491 326 0 3 22
0 13 9 14
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 1 0
1 U
9914 0 0
0
0
9 2-In XOR~
219 524 287 0 3 22
0 4 17 15
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 1 0
1 U
3747 0 0
0
0
9 2-In AND~
219 355 180 0 3 22
0 18 2 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
3549 0 0
0
0
12 Hex Display~
7 51 434 0 18 19
10 2 5 8 20 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
1 Y
-4 -38 3 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
7931 0 0
0
0
8 Hex Key~
166 87 502 0 11 12
0 8 2 2 2 0 0 0 0 0
0 48
0
0 0 4656 0
0
2 B3
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9325 0 0
0
0
8 Hex Key~
166 120 502 0 11 12
0 5 2 2 2 0 0 0 0 0
1 49
0
0 0 4656 0
0
2 B2
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8903 0 0
0
0
8 Hex Key~
166 153 501 0 11 12
0 2 2 2 2 0 0 0 0 0
0 48
0
0 0 4656 0
0
2 B1
-6 -35 8 -27
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3834 0 0
0
0
9 2-In XOR~
219 391 286 0 3 22
0 7 5 17
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 1 0
1 U
3363 0 0
0
0
9 Inverter~
13 207 184 0 2 22
0 19 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 2 0
1 U
7668 0 0
0
0
9 2-In XOR~
219 344 121 0 3 22
0 19 2 16
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 1446731082
65 0 0 0 4 1 1 0
1 U
4718 0 0
0
0
8 Hex Key~
166 67 232 0 11 12
0 3 3 3 3 0 0 0 0 0
0 48
0
0 0 4656 0
0
2 A3
-5 -34 9 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3874 0 0
0
0
8 Hex Key~
166 101 232 0 11 12
0 7 3 3 3 0 0 0 0 0
1 49
0
0 0 4656 0
0
2 A2
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6671 0 0
0
0
8 Hex Key~
166 134 232 0 11 12
0 19 3 3 3 0 0 0 0 0
1 49
0
0 0 4656 0
0
2 A1
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3789 0 0
0
0
12 Hex Display~
7 566 94 0 18 19
10 16 15 14 21 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
7 Resulta
-25 -38 24 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
4871 0 0
0
0
12 Hex Display~
7 23 125 0 18 19
10 19 7 3 22 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
1 X
-4 -38 3 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3750 0 0
0
0
7 Ground~
168 24 586 0 1 3
0 23
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
3 GND
8778 0 0
0
0
50
4 0 2 0 0 4096 0 13 0 0 27 2
144 525
144 580
3 0 2 0 0 0 0 13 0 0 27 2
150 525
150 580
2 0 2 0 0 0 0 13 0 0 27 2
156 525
156 580
4 0 2 0 0 0 0 11 0 0 27 2
78 526
78 580
3 0 2 0 0 0 0 11 0 0 27 2
84 526
84 580
2 0 2 0 0 0 0 11 0 0 27 2
90 526
90 580
4 0 3 0 0 4096 0 19 0 0 36 2
125 256
125 255
3 0 3 0 0 0 0 19 0 0 36 2
131 256
131 255
2 0 3 0 0 0 0 19 0 0 36 2
137 256
137 255
4 0 3 0 0 0 0 18 0 0 36 2
92 256
92 255
3 0 3 0 0 0 0 18 0 0 36 2
98 256
98 255
2 0 3 0 0 0 0 18 0 0 36 2
104 256
104 255
4 0 3 0 0 0 0 17 0 0 36 2
58 256
58 255
3 0 3 0 0 0 0 17 0 0 36 2
64 256
64 255
2 0 3 0 0 0 0 17 0 0 36 2
70 256
70 255
2 0 4 0 0 4224 0 3 0 0 19 5
536 515
299 515
299 433
438 433
438 427
1 0 5 0 0 4096 0 3 0 0 18 4
536 497
314 497
314 470
426 470
2 0 5 0 0 12416 0 4 0 0 30 4
536 478
426 478
426 470
198 470
2 0 4 0 0 128 0 5 0 0 42 5
536 435
536 427
428 427
428 195
436 195
1 0 6 0 0 4224 0 4 0 0 28 4
536 460
301 460
301 415
354 415
4 0 2 0 0 0 0 12 0 0 27 3
111 526
123 526
123 580
3 0 2 0 0 0 0 12 0 0 27 3
117 526
129 526
129 580
2 0 2 0 0 0 0 12 0 0 27 3
123 526
135 526
135 580
0 1 7 0 0 4096 0 0 6 49 0 4
363 282
275 282
275 353
283 353
0 3 8 0 0 8192 0 0 10 29 0 4
187 590
187 591
48 591
48 458
0 2 5 0 0 0 0 0 10 30 0 4
153 530
153 541
54 541
54 458
0 1 2 0 0 8192 0 0 10 46 0 4
192 525
192 580
60 580
60 458
1 2 6 0 0 128 0 5 6 0 0 4
536 417
354 417
354 353
319 353
1 2 8 0 0 12432 0 11 2 0 0 5
96 526
96 590
330 590
330 335
373 335
1 2 5 0 0 12416 0 12 14 0 0 6
129 526
129 530
198 530
198 298
375 298
375 295
4 2 9 0 0 4224 0 1 7 0 0 3
585 376
475 376
475 335
3 3 10 0 0 12416 0 3 1 0 0 5
581 506
581 515
463 515
463 385
539 385
3 2 11 0 0 8320 0 4 1 0 0 4
581 469
513 469
513 376
540 376
3 1 12 0 0 8320 0 5 1 0 0 5
581 426
581 434
376 434
376 367
539 367
3 1 13 0 0 8320 0 2 7 0 0 3
422 326
422 317
475 317
0 3 3 0 0 4096 0 0 21 37 0 3
150 255
20 255
20 149
1 1 3 0 0 16512 0 17 2 0 0 5
76 256
76 255
150 255
150 317
373 317
3 3 14 0 0 8320 0 7 20 0 0 3
524 326
563 326
563 118
3 2 15 0 0 4224 0 8 20 0 0 4
557 287
557 155
569 155
569 118
3 1 16 0 0 4224 0 16 20 0 0 3
377 121
575 121
575 118
3 2 17 0 0 4224 0 14 8 0 0 4
424 286
493 286
493 296
508 296
3 1 4 0 0 0 0 9 8 0 0 6
376 180
436 180
436 196
437 196
437 278
508 278
2 0 2 0 0 0 0 9 0 0 46 4
331 189
256 189
256 201
239 201
2 1 18 0 0 12416 0 15 9 0 0 4
228 184
243 184
243 171
331 171
0 1 19 0 0 8192 0 0 15 50 0 3
212 158
192 158
192 184
1 2 2 0 0 8320 0 13 16 0 0 4
162 525
239 525
239 130
328 130
0 2 7 0 0 8192 0 0 21 49 0 4
168 277
168 170
26 170
26 149
0 1 19 0 0 8192 0 0 21 50 0 4
158 158
158 179
32 179
32 149
1 1 7 0 0 8320 0 18 14 0 0 7
110 256
110 277
363 277
363 282
363 282
363 277
375 277
1 1 19 0 0 16512 0 19 16 0 0 7
143 256
143 250
158 250
158 158
324 158
324 112
328 112
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3999480 1079360 100 100 0 0
0 0 0 0
1 66 162 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
